//apb defines file
`define uvm_apb_dsize 32
`define uvm_apb_asize 32
