//i2s_uvc interface
//author: astrakhov, JSC MERI
//date: 31.10.2021

interface i2s_uvc_interface (
  input logic TCLK
);

logic WS;
logic TD;

endinterface
