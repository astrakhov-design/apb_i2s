//i2s uvm package
//author: astrakhov, JSC MERI
//date: 05.11.2021
package i2s_pkg;
  import uvm_pkg::*;
  `include "i2s_seq_item.svh"
  `include "i2s_seq_lib.svh"
  `include "i2s_monitor.svh"
  `include "i2s_agent.svh"
  `include "i2s_scb.svh"
  `include "i2s_env.svh"

endpackage
