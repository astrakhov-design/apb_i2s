//register address definition list
`define CR_ADDR   32'h00
`define SR_ADDR   32'h04
`define TXR_ADDR  32'h08
`define TXL_ADDR  32'h0C
