package apb_pkg;
  import uvm_pkg::*;
  `include "apb_defines.svh"
  `include "apb_seq_item.svh"
  `include "apb_sequencer.svh"
  `include "apb_seq_lib.svh"
  `include "apb_driver.svh"
  `include "apb_monitor.svh"
  `include "apb_agent.svh"
  `include "apb_scb.svh"
  `include "apb_env.svh"

endpackage
